$SRLatch [
	s*;
	r*;
	q: nor s p;
	p: nor r q;
]

sr#SRLatch*;
i1: hi;
i2: lo;
sr.s: i1;
sr.r: i2;